`ifndef __WIDTHS_VH
`define __WIDTHS_VH 1

`define LEN_W 10
`define TD_W 1

`define BARDECODE_W 8
`define OFFSET_W 4
`define EP_W 1
`define TC_W 3
`define TYPE_W 5
`define ATTR_W 3
`define FMT_W 3
`define FBE_W 4
`define LBE_W 4
`define TAG_W 8
`define ADDR_W 64
`define REQID_W 16
`define CPLID_W 16
`define BYTECNT_W 12
`define STAT_W 3
`define LOWADDR_W 7

`define EXT_TYPE_W 3

`define LINKWIDTH_W 6
`define LINKRATE_W 4
`define MAXREAD_W 3
`define MAXPAYLOAD_W 3

`define PCIE_CONFIGURATION_REGISTER_WIDTH 16
`define PCIE_BUS_ID_WIDTH 8
`define PCIE_DEVICE_ID_WIDTH 5
`define PCIE_FUNCTION_ID_WIDTH 3

`endif

